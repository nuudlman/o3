
module o3_top
(
    input bit clk,
    input bit rst
);

    initial
    begin
        $finish();
    end

endmodule